// There is nothing here, really.
