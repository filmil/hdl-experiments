-- The library here is ex4_lib1.

--! @package lib1
--! @brief A library package containing a simple constant.
package lib1 is
    
   -- This is ex4_lib1.lib1.c
   --! @constant c
   --! @brief An integer constant initialized to 1.
   constant c: integer := 1; 
    
end package lib1;
